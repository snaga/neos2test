module main(input clk, input reset);

    main u0 (
		.clk_clk (clk),
		.reset_reset_n (reset)
	 );

endmodule
